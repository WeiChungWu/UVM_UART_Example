`include "uart_ip_tb.sv"
`include "uart_base_test.sv"
`include "uart_rdwr_test.sv"
